module NIOS_proj ();





endmodule 