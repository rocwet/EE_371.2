
module first_nios2_system (
	clk_clk,
	reset_reset_n,
	led_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	led_connection_export;
endmodule
